module tb();
  logic [3:0]a;
  logic y;
  XOR_4 dut([3:0]a,y);

initial begin
  $dumpfile("dump.vcd");
	$dumpvars;
  a[0]=0;a[1]=0;a[2]=0;a[3]=0;
  #10 a[0]=0;a[1]=0;a[2]=0;a[3]=1;
  #10 a[0]=0;a[1]=0;a[2]=1;a[3]=0;
  #10 a[0]=0;a[1]=0;a[2]=1;a[3]=1;
  #10 a[0]=0;a[1]=1;a[2]=0;a[3]=0;
  #10 a[0]=0;a[1]=1;a[2]=0;a[3]=1;
  #10 a[0]=0;a[1]=1;a[2]=1;a[3]=0;
  #10 a[0]=0;a[1]=1;a[2]=1;a[3]=1;
  #10 a[0]=1;a[1]=0;a[2]=0;a[3]=0;
  #10 a[0]=1;a[1]=0;a[2]=0;a[3]=1;
  #10 a[0]=1;a[1]=0;a[2]=1;a[3]=0;
  #10 a[0]=1;a[1]=0;a[2]=1;a[3]=1;
  #10 a[0]=1;a[1]=1;a[2]=0;a[3]=0;
  #10 a[0]=1;a[1]=1;a[2]=0;a[3]=1;
  #10 a[0]=1;a[1]=1;a[2]=1;a[3]=0;
  #10 a[0]=1;a[1]=1;a[2]=1;a[3]=1;
end
endmodule

  
